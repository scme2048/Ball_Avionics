//////////////////////////////////////////////////////////////////////
// Created by Microsemi SmartDesign Tue Jan 12 11:57:26 2016
// Testbench Template
// This is a basic testbench that instantiates your design with basic 
// clock and reset pins connected.  If your design has special
// clock/reset or testbench driver requirements then you should 
// copy this file and modify it. 
//////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: timestamp_testbench.v
// File history:
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// <Description here>
//
// Targeted device: <Family::ProASIC3L> <Die::A3PE3000L> <Package::484 FBGA>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

`timescale 1ns/100ps

module timestamp_testbench;

parameter SYSCLK_PERIOD = 100000000;// 10HZ

reg SYSCLK;
reg NSYSRESET;

initial
begin
    SYSCLK = 1'b0;
    NSYSRESET = 1'b0;
end

//////////////////////////////////////////////////////////////////////
// Reset Pulse
//////////////////////////////////////////////////////////////////////
initial
begin
    #(SYSCLK_PERIOD * 10 )
        NSYSRESET = 1'b1;
end


//////////////////////////////////////////////////////////////////////
// Clock Driver
//////////////////////////////////////////////////////////////////////
always @(SYSCLK)
    #(SYSCLK_PERIOD / 2.0) SYSCLK <= !SYSCLK;

wire [23:0] ts_out;
//////////////////////////////////////////////////////////////////////
// Instantiate Unit Under Test:  timestamp
//////////////////////////////////////////////////////////////////////
timestamp timestamp_0 (
    // Inputs
    .CLK_10HZ(SYSCLK),
    .RESET(NSYSRESET),

    // Outputs
    .TIMESTAMP( ts_out)

    // Inouts

);

endmodule

