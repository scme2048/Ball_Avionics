///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: spi_interface.v
//
// Description: 
// Transceiver interface. Commands mode for tx/rx as well as data tx/rx.
//
// <Description here>
//
// Targeted device: <Family::ProASIC3L> <Die::A3PE3000L> <Package::484 FBGA>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

//`timescale <time_units> / <precision>

module spi_interface( port1, port2, port3, port4 );
input port1, port2;
output port3;
inout port4;

//<statements>

endmodule

