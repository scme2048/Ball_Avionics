///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: write_address_traversal.v
// File history:
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// <Description here>
//
// Targeted device: <Family::ProASIC3L> <Die::A3PE3000L> <Package::484 FBGA>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

//`timescale <time_units> / <precision>

module write_address_traversal( port1, port2, port3, port4 );
input port1, port2;
output port3;
inout port4;

//<statements>

endmodule

